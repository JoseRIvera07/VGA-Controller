module sprite(
	input clk,
	input [3:0] step,
	input [2:0] cuadrante,
	input [9:0] pixel_x,pixel_y,
	output enable,
	output logic [4:0] sprite
);
/*
COLORES
[
'0x00000000', 00000, 000000000000000000000000
'0xff582818', 00001, 101100001010000011000000
'0xff784820', 00010, 111100001001000010000000
'0xffe8e0e0', 00011, 111010001110000011100000
'0xff381810', 00100, 111000001100000010000000
'0xff181818', 00101, 110000001100000011000000
'0xff203068', 00110, 100000001100000011010000
'0xfff8f8f8', 00111, 111110001111100011111000
'0xff4078d8', 01000, 100000001111000011011000
'0xff80b0f8', 01001, 100000001011000011111000
'0xff1810c0', 01010, 110000001000000011000000
'0xff6848e8', 01011, 110100001001000011101000
'0xff9878e8', 01100, 100110001111000011101000
'0xff5020c8', 01101, 101000001000000011001000
'0xff505048', 01110, 101000001010000010010000
'0xff103868', 01111, 100000001110000011010000
'0xffa8b090', 10000, 101010001011000010010000
'0xff206090', 10001, 100000001100000010010000
'0xff102048', 10010, 100000001000000010010000
'0xffa0f8f8', 10011, 101000001111100011111000
'0xff000000', 10100, 000000000000000000000000
'0xff48e0f0', 10101, 100100001110000011110000
'0xff181068', 10110, 110000001000000011010000
'0xff1038f8'  10111, 100000001110000011111000
]
*/

logic [0:4]RAM [0:63] [0:63]  = '{
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00001, 5'b00001, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00001, 5'b00001, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00001, 5'b00001, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00010, 5'b00010, 5'b00100, 5'b00100, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00001, 5'b00001, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00010, 5'b00010, 5'b00100, 5'b00100, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00100, 5'b00100, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00001, 5'b00001, 5'b00100, 5'b00100, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00100, 5'b00100, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00001, 5'b00001, 5'b00100, 5'b00100, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00001, 5'b00001, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00001, 5'b00001, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00100, 5'b00100, 5'b00001, 5'b00001, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00001, 5'b00001, 5'b00100, 5'b00100, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00100, 5'b00100, 5'b00001, 5'b00001, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00001, 5'b00001, 5'b00100, 5'b00100, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00100, 5'b00100, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00100, 5'b00100, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00101, 5'b00101, 5'b00110, 5'b00110, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00101, 5'b00101, 5'b00110, 5'b00110, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00101, 5'b00101, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b01000, 5'b01000, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00111, 5'b00111, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00101, 5'b00101, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b01000, 5'b01000, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00111, 5'b00111, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00110, 5'b00110, 5'b01000, 5'b01000, 5'b01001, 5'b01001, 5'b00110, 5'b00110, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b01010, 5'b01010, 5'b00111, 5'b00111, 5'b01001, 5'b01001, 5'b00111, 5'b00111, 5'b01010, 5'b01010, 5'b00111, 5'b00111, 5'b00110, 5'b00110, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00110, 5'b00110, 5'b01000, 5'b01000, 5'b01001, 5'b01001, 5'b00110, 5'b00110, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b01010, 5'b01010, 5'b00111, 5'b00111, 5'b01001, 5'b01001, 5'b00111, 5'b00111, 5'b01010, 5'b01010, 5'b00111, 5'b00111, 5'b00110, 5'b00110, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00110, 5'b00110, 5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b00101, 5'b00101, 5'b01001, 5'b01001, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01101, 5'b01101, 5'b00110, 5'b00110, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00110, 5'b00110, 5'b01000, 5'b01000, 5'b01000, 5'b01000, 5'b00101, 5'b00101, 5'b01001, 5'b01001, 5'b00111, 5'b00111, 5'b00111, 5'b00111, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01100, 5'b01100, 5'b01100, 5'b01100, 5'b01101, 5'b01101, 5'b00110, 5'b00110, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b01000, 5'b01000, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b01001, 5'b01001, 5'b01011, 5'b01011, 5'b01101, 5'b01101, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01100, 5'b01100, 5'b01101, 5'b01101, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b01000, 5'b01000, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b01001, 5'b01001, 5'b01011, 5'b01011, 5'b01101, 5'b01101, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01011, 5'b01100, 5'b01100, 5'b01101, 5'b01101, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b01000, 5'b01000, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b01000, 5'b01000, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b01101, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b01000, 5'b01000, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b00110, 5'b00110, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b00110, 5'b00110, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b01000, 5'b01000, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b00110, 5'b00110, 5'b01001, 5'b01001, 5'b01001, 5'b01001, 5'b00110, 5'b00110, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b00000, 5'b00000, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00100, 5'b00100, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00100, 5'b00100, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b00000, 5'b00000, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00100, 5'b00100, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00100, 5'b00100, 5'b00110, 5'b00110, 5'b00110, 5'b00110, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b01110, 5'b01110, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b01110, 5'b01110, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b01111, 5'b01111, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00010, 5'b00010, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00101, 5'b00101, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b01110, 5'b01110, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b01110, 5'b01110, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b01111, 5'b01111, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00010, 5'b00010, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00101, 5'b00101, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b10000, 5'b10000, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b01110, 5'b01110, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b01111, 5'b01111, 5'b10001, 5'b10001, 5'b00001, 5'b00001, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00100, 5'b00100, 5'b00101, 5'b00101, 5'b01110, 5'b01110, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b10000, 5'b10000, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b01110, 5'b01110, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b01111, 5'b01111, 5'b10001, 5'b10001, 5'b00001, 5'b00001, 5'b00010, 5'b00010, 5'b00010, 5'b00010, 5'b00100, 5'b00100, 5'b00101, 5'b00101, 5'b01110, 5'b01110, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b10000, 5'b10000, 5'b00101, 5'b00101, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b01111, 5'b01111, 5'b10001, 5'b10001, 5'b00001, 5'b00001, 5'b00010, 5'b00010, 5'b00100, 5'b00100, 5'b00101, 5'b00101, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b00011, 5'b00011, 5'b00011, 5'b00011, 5'b10000, 5'b10000, 5'b00101, 5'b00101, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b01111, 5'b01111, 5'b10001, 5'b10001, 5'b00001, 5'b00001, 5'b00010, 5'b00010, 5'b00100, 5'b00100, 5'b00101, 5'b00101, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00001, 5'b00001, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00101, 5'b00101, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b10000, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00001, 5'b00001, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b00001, 5'b00001, 5'b00001, 5'b00001, 5'b00100, 5'b00100, 5'b00100, 5'b00100, 5'b00101, 5'b00101, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b01110, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b10001, 5'b10001, 5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10011, 5'b10011, 5'b10010, 5'b10010, 5'b10100, 5'b10100, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b10001, 5'b10001, 5'b10011, 5'b10011, 5'b10011, 5'b10011, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10011, 5'b10011, 5'b10010, 5'b10010, 5'b10100, 5'b10100, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b01111, 5'b01111, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10101, 5'b10101, 5'b10110, 5'b10110, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b01111, 5'b01111, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10101, 5'b10101, 5'b10101, 5'b10101, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10101, 5'b10101, 5'b10110, 5'b10110, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b10010, 5'b10010, 5'b01111, 5'b01111, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10010, 5'b10010, 5'b01111, 5'b01111, 5'b10110, 5'b10110, 5'b10111, 5'b10111, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b10010, 5'b10010, 5'b01111, 5'b01111, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10010, 5'b10010, 5'b01111, 5'b01111, 5'b10110, 5'b10110, 5'b10111, 5'b10111, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01111, 5'b01111, 5'b00101, 5'b00101, 5'b10010, 5'b10010, 5'b01111, 5'b01111, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b01111, 5'b01111, 5'b10010, 5'b10010, 5'b10111, 5'b10111, 5'b01010, 5'b01010, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b01111, 5'b01111, 5'b00101, 5'b00101, 5'b10010, 5'b10010, 5'b01111, 5'b01111, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b01111, 5'b01111, 5'b10010, 5'b10010, 5'b10111, 5'b10111, 5'b01010, 5'b01010, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b01010, 5'b01010, 5'b10110, 5'b10110, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b01111, 5'b01111, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b01111, 5'b01111, 5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b01010, 5'b01010, 5'b10110, 5'b10110, 5'b01111, 5'b01111, 5'b01111, 5'b01111, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b01111, 5'b01111, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b10001, 5'b01111, 5'b01111, 5'b01010, 5'b01010, 5'b01010, 5'b01010, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b01111, 5'b01111, 5'b10001, 5'b10001, 5'b01010, 5'b01010, 5'b10110, 5'b10110, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b10010, 5'b10010, 5'b10010, 5'b10010, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b01111, 5'b01111, 5'b10001, 5'b10001, 5'b01010, 5'b01010, 5'b10110, 5'b10110, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b10110, 5'b10110, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b10110, 5'b10110, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b10110, 5'b10110, 5'b10110, 5'b10110, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00101, 5'b00101, 5'b00101, 5'b00101, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000},
 '{5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000, 5'b00000}
 };
 

always @(posedge clk)
begin
	if(step==4'b0010)
	begin
		if(cuadrante==3'b001)
		begin
			if(pixel_x>=266 && pixel_x < 330 && pixel_y>= 120 && pixel_y < 184)
			begin
				sprite <= RAM[pixel_y-120][pixel_x-266];
				enable <= 1;
			end
			else begin
				enable <= 0;
			end
		end

		else if(cuadrante==3'b010)
		begin
			if(pixel_x>=586 && pixel_x < 650 && pixel_y>= 120 && pixel_y < 184)
			begin
				sprite <= RAM[pixel_y-120][pixel_x-586];
				enable <= 1;
			end
			else begin
				enable <= 0;
			end
		end
		
		else if(cuadrante==3'b011)
		begin
			if(pixel_x>=266 && pixel_x < 330 && pixel_y>= 361 && pixel_y < 425)
			begin
				sprite <= RAM[pixel_y-361][pixel_x-266];
				enable <= 1;
			end
			else begin
				enable <= 0;
			end
		end
		
		else if(cuadrante==3'b100)
		begin
			if(pixel_x>=586 && pixel_x < 650 && pixel_y>= 361 && pixel_y < 425)
			begin
				sprite <= RAM[pixel_y-361][pixel_x-586];
				enable <= 1;
			end
			else begin
				enable <= 0;
			end
		end
		else enable <= 0;
	end
	else enable <= 0;

end
endmodule
